module and_module (
    in_1, // input
    in_2, // input
    out   // output
);

    input in_1;
    input in_2;
    output out;

    assign out = in_1 && in_2;
    
endmodule
